
module Problema_3_tb;

  // Parameters
  parameter N = 4;

  // Inputs for substractor
  logic a, b, c_in;

  // Outputs for substractor
  logic result, c_out;

  // Inputs for Problema_3
  logic [N-1:0] a_vec, b_vec;

  // Outputs for Problema_3
  logic [N-1:0] result_vec;
  logic neg_flag, zr_flag, cry_flag, of_flag;

  // Instantiate the substractor module
  substractor uut_substractor (
    .a(a),
    .b(b),
    .c_in(c_in),
    .result(result),
    .c_out(c_out)
  );

  // Instantiate the Problema_3 module
  Problema_3 #(.N(N)) uut_Problema_3 (
    .a(a_vec),
    .b(b_vec),
    .result(result_vec),
    .neg_flag(neg_flag),
    .zr_flag(zr_flag),
    .cry_flag(cry_flag),
    .of_flag(of_flag)
  );

  initial begin
    // Test Case 1: 0 - 0 - 0 = 0, No carry
    a = 0; b = 0; c_in = 0;
    #30;

    // Test Case 2: 0 - 1 - 0 = 1, Carry generated
    a = 0; b = 1; c_in = 0;
    #30;

    // Test Case 3: 1 - 1 - 1 = 1, Carry generated
    a = 1; b = 1; c_in = 1;
    #30;

    // Test Case 4: 1 - 0 - 1 = 0, No carry
    a = 1; b = 0; c_in = 1;
    #30;
  end

  initial begin
    
    // Test Case 1: 4'b0000 - 4'b0000 = 4'b0000
    a_vec = 4'b0000; b_vec = 4'b0000;
    #30;

    // Test Case 2: 4'b0001 - 4'b0001 = 4'b0000
    a_vec = 4'b0001; b_vec = 4'b0001;
    #30;

    // Test Case 3: 4'b1111 - 4'b0001 = 4'b1110
    a_vec = 4'b1111; b_vec = 4'b0001;
    #30;

    // Test Case 4: 4'b0111 - 4'b1000 = 4'b1111
    a_vec = 4'b0111; b_vec = 4'b1000;
    #30;

    // Test Case 5: 4'b1000 - 4'b1000 = 4'b0000
    a_vec = 4'b1000; b_vec = 4'b1000;
    #30;
	 
    // Test Case 6: 4'b1010 - 4'b0101 = 4'b0101
    a_vec = 4'b1010; b_vec = 4'b0101;
    #30;

    // Test Case 7: 4'b0011 - 4'b0110 = 4'b1101
    a_vec = 4'b0011; b_vec = 4'b0110;
    #30;
  end

endmodule
